library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;
library cplxlib;
  use cplxlib.cplx_pkg.all;
library dsplib;

-- Version V2 - uses cplx_mult_accu
-- INPUT  = row vector (stream of single input values)
-- OUTPUT = column vector (all output values parallel in one cycle)

entity dft8_v2 is
port (
  clk      : in  std_logic; -- clock
  rst      : in  std_logic; -- reset
  inverse  : in  std_logic := '0'; -- inverse FFT
  start    : in  std_logic; -- start pulse
  idx_in   : in  unsigned(2 downto 0);
  data_in  : in  cplx;
  data_out : out cplx_vector(0 to 7) := cplx_vector_reset(18,8,"R")
);
end entity;

-------------------------------------------------------------------------------

architecture rtl of dft8_v2 is

  constant DFTMTX_RESOLUTION : positive range 8 to 32 := 16; -- Real/Imag width in bits
  constant DFTMTX_POWER_LD : positive := DFTMTX_RESOLUTION-1;

  signal fft_start : std_logic := '0';
  signal fft_in : cplx := cplx_reset(18,"R");

  signal dftmtx_slv : std_logic_vector(8*2*DFTMTX_RESOLUTION-1 downto 0);
  signal dftmtx_16bit : cplx16_vector(0 to 7);
  signal dftmtx_18bit : cplx_vector(0 to 7);

  signal run : std_logic := '0';
  signal inverse_q,conj : std_logic := '0';
  signal idx : unsigned(2 downto 0);

  constant MAX_NUM_PIPE_DSP : positive := 10;
  
  type natural_vector is array(integer range <>) of natural;
  signal PIPESTAGES : natural_vector(0 to 7);

  type t_idx is array(integer range <>) of unsigned(2 downto 0);
  signal idx_q : t_idx(0 to MAX_NUM_PIPE_DSP);

  signal data_out_i : cplx_vector(0 to 7);

begin

  -- data input
  p_din : process(clk)
  begin
    if rising_edge(clk) then
      if start='1' or run='0' then
        inverse_q <= inverse;
      end if;
      fft_in <= data_in;
      fft_start <= start;
    end if;
  end process;

  -- input index generation
  p_idx : process(clk)
  begin
    if rising_edge(clk) then
      if rst='1' then
        idx <= (others=>'0');
        run <= '0';

      elsif (start='1' or run='1') then
        if data_in.vld='1' then
          if idx=7 then
            idx <= (others=>'0');
            run <= '0';
          else
            idx <= idx + 1;
            run <= '1';
          end if;
        end if;
      else
        idx <= (others=>'0');
        run <= '0';
     end if; --reset
    end if; --clock
  end process;

  conj <= inverse when start='1' else inverse_q;

  -- DFT-Matrix ROM,  one cycle delay
  i_dtfmtx : entity work.dftmtx8
  generic map(
    IQ_WIDTH => DFTMTX_RESOLUTION,
    POWER_LD => DFTMTX_POWER_LD
  )
  port map(
    clk  => clk,
    rst  => rst,
    idx  => idx,
    conj => conj,
    dout => dftmtx_slv
  );

  -- ROM output data to complex vector
  dftmtx_16bit <= to_cplx_vector(slv=>dftmtx_slv, n=>8, vld=>'1');
  dftmtx_18bit <= resize(dftmtx_16bit,18); -- resize to 18-bit standard for VHDL-1993

  g_loop : for n in 0 to 7 generate
  -- multiplier
  i_mult : entity cplxlib.cplx_mult_accu
  generic map(
    NUM_MULT => 1,
    NUM_SUMMAND => 8,
    NUM_INPUT_REG => 1,
    NUM_OUTPUT_REG => 0,
    OUTPUT_SHIFT_RIGHT => DFTMTX_POWER_LD,
    MODE => "NSO" -- round + saturation + overflow detection
  )
  port map(
    clk        => clk,
    clk2       => open, -- unused
    clr        => fft_start,
    neg        => "0",
    x(0)       => fft_in,
    y(0)       => dftmtx_18bit(n),
    result     => data_out_i(n),
    PIPESTAGES => PIPESTAGES(n)
  );
  end generate;

  -- bypassed index
  idx_q(0) <= idx;
  g_delay : for n in 1 to MAX_NUM_PIPE_DSP generate
    idx_q(n) <= idx_q(n-1) when rising_edge(clk);
  end generate;

  p_out : process(clk)
  begin
    if rising_edge(clk) then
      if idx_q(PIPESTAGES(0)+1)=7 then
        data_out <= data_out_i;
      else
        for n in 0 to 7 loop
          data_out(n).vld <= '0';
        end loop;
      end if;
    end if;
  end process;

end architecture;
